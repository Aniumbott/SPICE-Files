* DC analysis of a NMOS transistor
.include "../Dependencies/cmos_90nm.txt"
M1 d g 0 0 NMOS w=0.25u L=0.9u
Vds d 0 1.2
Vgs g 0 1.2

* DC analysis
.dc Vds 0.1 1.2 0.001

.control
run
set color0 = white;
set xbrushwidth = 3.5;
plot -i(Vds) 
.endc
.end