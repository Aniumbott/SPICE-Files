* *Transient Analysis of TTL Inverter
.MODEL bjt npn(BF=20)
Q1 c1 b1 e1 bjt
Q2 c2 c1 0 bjt
Rb b1 cc 10k
Rc c2 cc 1k
Vcc cc 0 5
Vin e1 0 5

* Transient analysis
.tran 0.1ps 40ns

.control 
run 
set color0=white
set xbrushwidth = 3
plot v(c2) v(e1) 
.endc
.end
