*Forward biased diode characteristics
.model mode1 d(n=2 Is=1E-12 Rs=10 Cjo=5p Tt=10n Vj=1 Bv=10)
vin 1 0 dc 5 
d1 2 0 mode1
r1 1 2 6.5k

*simulation
.dc vin 0 5 0.05

.control
run
set color0=white
set xbrushwidth=3.5
plot -i (vin)
.endc
.end
