*pmos u20ec055
.include cmos_130nm.txt
M1 D G S Su PMOS W=1u L=0.13u
Vs  S 0 0v
Vsu Su 0 0v
Vgs G S 1.2v
Vds D S -1.2V
.dc Vgs -2 0 0.01
*.dc Vds -1.2 0 0.01
.control
run
plot i(Vds)
.endc
.end