* Fanout of TTL 
.MODEL bjt npn(BF=20)

* Subcircuit for TTL inverter
.subckt ttl_inv in cc out
    Rb b1 cc 10k
    Rc out cc 1k
    Q1 c1 b1 in bjt
    Q2 out c1 0 bjt
.ends ttl_inv

Vcc cc 0 5
Vin in 0 5

* Fanout 
xmaster in cc out ttl_inv

x1 out cc out1 ttl_inv
x2 out cc out2 ttl_inv
x3 out cc out3 ttl_inv
x4 out cc out4 ttl_inv
x5 out cc out5 ttl_inv
x6 out cc out6 ttl_inv
x7 out cc out7 ttl_inv
x8 out cc out8 ttl_inv
x9 out cc out9 ttl_inv
x10 out cc out10 ttl_inv
x11 out cc out11 ttl_inv
x12 out cc out12 ttl_inv

* VTC using DC analysis
.dc Vin 0 5 0.1

.control 
run 
set color0=white
set xbrushwidth = 3
plot v(in) v(out) 
.endc
.end
