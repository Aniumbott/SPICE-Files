*Fanout of RTL 
.model bjt npn (Bf=20)

Q1 2 1 0 bjt
Rb 4 1 10k
Rc 2 3 1k
Vcc 3 0 5
Vin 4 0 5

* Subcircuit of RTL
.subckt rtl out in c 0
Q2 out y 0 bjt
Rb1 in y 10k
Rc1 c out 1k
.ends rtl

x1 out1 2 3 0 rtl
x2 out2 2 3 0 rtl
x3 out3 2 3 0 rtl
x4 out4 2 3 0 rtl
x5 out5 2 3 0 rtl
x6 out6 2 3 0 rtl
x7 out7 2 3 0 rtl

* DC analysis
.dc Vin 0 5 0.05

.control
run
set color0=white
set xbrushwidth=3.5
plot V(2) V(4)
.endc
.end
