*Voltage Transfer Characteristics (VTC) and Noise Margin (NM) of RTL inverter
.model bjt NPN (BF=20)

Q1 2 1 0 bjt
Rc 2 3 1k
Rb 4 1 10k
Vcc 3 0 5
Vin 4 0 5

* VTC using DC analysis
.dc Vin 0 5 0.05

.control
run
set color0=white
set xbrushwidth=3.5
plot v(2) 
plot v(4)
plot v(2) v(4)
.endc
.end
