*Transient Analysis of RTL Inverter
.model bjt NPN (BF=20)

Q 2 1 0 bjt
Rc 2 3 1k
Rb 4 1 10k
Vcc 3 0 5
Vin 4 0 pulse (0 5 1ns 1ns 11ns 40us 80us)
c1 2 0 1p

* Transient Analysis
.tran 1ns 160us

.control
run
set color0=white
set xbrushwidth=3.5
plot v(4) 
plot v(2)
plot v(4) v(2)
.endc 
.end
